module e;
	always #1 $write("e");
endmodule